//--------------------------------------------------------------
/*
    Filename: core.v

    RV32I top module.
*/
//--------------------------------------------------------------

module core (

);



endmodule : core