//--------------------------------------------------------------
/*
    Filename: D_stage.v

    Decode stage top module.
*/
//--------------------------------------------------------------

module D_stage (

);



endmodule : D_stage