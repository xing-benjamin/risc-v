//--------------------------------------------------------------
/*
    Filename: M_stage.v

    Memory stage top module.
*/
//--------------------------------------------------------------

module M_stage (

);



endmodule : M_stage