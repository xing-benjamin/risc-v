//--------------------------------------------------------------
/*  
    Filename: dl_xor.v

    Paramterized bitwise XOR operation.
*/
//--------------------------------------------------------------

`ifndef __DL_XOR_V__
`define __DL_XOR_V__

module dl_xor #(
    parameter   NUM_BITS = 1
)(
    // TODO EMILY: define input and output ports
);
    // TODO EMILY: implement bitwise XOR

endmodule

`endif // __DL_XOR_V__