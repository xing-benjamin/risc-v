//--------------------------------------------------------------
/*  
    Filename: dl_or.v

    Paramterized bitwise OR operation.
*/
//--------------------------------------------------------------

`ifndef __DL_OR_V__
`define __DL_OR_V__

module dl_or #(
    parameter   NUM_BITS = 1
)(
    // TODO EMILY: define input and output ports
);
    // TODO EMILY: implement bitwise OR

endmodule

`endif // __DL_OR_V__