//--------------------------------------------------------------
/*  
    Filename: dl_and.v

    Paramterized bitwise AND operation.
*/
//--------------------------------------------------------------

`ifndef __DL_AND_V__
`define __DL_AND_V__

module dl_and #(
    parameter   NUM_BITS = 1
)(
    // TODO EMILY: define input and output ports
);
    // TODO EMILY: implement bitwise AND

endmodule

`endif // __DL_AND_V__