//--------------------------------------------------------------
/*
    Filename: F_stage.v

    Fetch stage top module.
*/
//--------------------------------------------------------------

module F_stage (

);



endmodule : F_stage