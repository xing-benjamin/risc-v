//--------------------------------------------------------------
/*
    Filename: W_stage.v

    Write stage top module.
*/
//--------------------------------------------------------------

module W_stage (

);



endmodule : W_stage